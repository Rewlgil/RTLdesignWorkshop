module remme (clk, reset, r, m);

  input clk, reset;
  input [3:0] r;
  output [3:0] m;




endmodule
