module vend (clk, reset, a, b, t, c);
  input clk, reset, a, b;
  output t, c;




endmodule
