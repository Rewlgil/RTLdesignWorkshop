module signed2twos (s, t);
  input [7:0] s;
  output [7:0] t;



endmodule
