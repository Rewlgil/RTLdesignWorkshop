module arb (clk, reset, req_a, req_b, grant_a, grant_b);

  input clk, reset;
  input req_a, req_b;
  output grant_a, grant_b;





endmodule
