module flt (clk, reset, n, t, n_best, t_best);
  input clk, reset;
  input [1:0] n;
  input [7:0] t;
  output [1:0] n_best;
  output [7:0] t_best;




endmodule
