module crossbar (in0, in1, in2, select, out0, out1, out2, valid);
  input [7:0] in0, in1, in2;
  input [5:0] select;
  output [7:0] out0, out1, out2;
  output valid;







endmodule
