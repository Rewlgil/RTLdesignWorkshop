module majority (a, b, c, m);
  input a, b, c;
  output m;

endmodule
