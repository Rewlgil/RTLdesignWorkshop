module signed_mag_compare (a, b, aLTb, aGTb, aEQb);
        
  input [6:0] a, b;
  output aLTb, aGTb, aEQb;








endmodule
